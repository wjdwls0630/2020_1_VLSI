** Generated for: hspiceD
** Generated on: Apr 18 15:53:12 2020
** Design library name: Library_Jin
** Design cell name: and2
** Design view name: schematic



** Library name: Library_Jin
** Cell name: nand2
** View name: schematic
.subckt nand2 a b gnd vdd y
m1 y b vdd vdd PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m0 y a vdd vdd PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m2 y a n1 gnd NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m3 n1 b gnd gnd NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
.ends nand2
** End of subcircuit definition.

** Library name: Library_Jin
** Cell name: inverter
** View name: schematic
.subckt inverter gnd input output vdd
m0 output input gnd gnd NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m1 output input vdd vdd PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
.ends inverter
** End of subcircuit definition.

** Library name: Library_Jin
** Cell name: and2
** View name: schematic
.subckt and2 y a b vdd gnd 
xi0 a b gnd vdd net10 nand2
xi1 gnd net10 y vdd inverter
.ends and2
