* SPICE NETLIST
***************************************

.SUBCKT TGFA_2010 B VDD A GND Cout Cin Sum
** N=12 EP=7 IP=0 FDC=14
M0 12 A 4 GND NMOS_VTL L=5e-08 W=9e-08 AD=2.655e-14 AS=1.62e-14 PD=7.7e-07 PS=5.4e-07 $X=-13995 $Y=4260 $D=1
M1 GND B 12 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.755e-14 AS=2.655e-14 PD=5.7e-07 PS=7.7e-07 $X=-13305 $Y=4260 $D=1
M2 Cout 5 A GND NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6875e-14 PD=5.45e-07 PS=5.55e-07 $X=-13270 $Y=3575 $D=1
M3 Sum 5 Cin GND NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6875e-14 PD=5.45e-07 PS=5.55e-07 $X=-12085 $Y=3570 $D=1
M4 5 4 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.125e-14 AS=1.1025e-14 PD=4.3e-07 PS=4.25e-07 $X=-11620 $Y=4290 $D=1
M5 Cout 4 Cin GND NMOS_VTL L=5e-08 W=9e-08 AD=1.665e-14 AS=1.665e-14 PD=5.5e-07 PS=5.5e-07 $X=-10755 $Y=3570 $D=1
M6 Sum Cin 5 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6425e-14 PD=5.45e-07 PS=5.45e-07 $X=-10625 $Y=4280 $D=1
M7 4 A B VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=5.31e-14 AS=3.195e-14 PD=9.5e-07 PS=7.15e-07 $X=-13995 $Y=5790 $D=0
M8 A B 4 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.51e-14 AS=5.31e-14 PD=7.5e-07 PS=9.5e-07 $X=-13305 $Y=5790 $D=0
M9 Cout 4 A VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.375e-14 PD=7.05e-07 PS=7.35e-07 $X=-13260 $Y=1815 $D=0
M10 Sum 4 Cin VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.195e-14 AS=3.465e-14 PD=7.15e-07 PS=7.45e-07 $X=-12075 $Y=1810 $D=0
M11 5 4 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.205e-14 AS=2.16e-14 PD=6.05e-07 PS=6e-07 $X=-11620 $Y=5790 $D=0
M12 Cout 5 Cin VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.375e-14 PD=7.05e-07 PS=7.35e-07 $X=-10740 $Y=1810 $D=0
M13 Sum Cin 4 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.465e-14 AS=3.06e-14 PD=7.45e-07 PS=7e-07 $X=-10625 $Y=5790 $D=0
.ENDS
***************************************
