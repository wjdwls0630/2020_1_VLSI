* SPICE NETLIST
***************************************

.SUBCKT NTAP_CDNS_592557639821
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PTAP_CDNS_592557639820
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pass_mux GND VDD C B A OUT
** N=6 EP=6 IP=2 FDC=2
M0 OUT C B GND NMOS_VTL L=5e-08 W=1.775e-07 AD=2.75125e-14 AS=2.6625e-14 PD=6.65e-07 PS=6.55e-07 $X=-13305 $Y=9245 $D=1
M1 OUT C A VDD PMOS_VTL L=5e-08 W=1.775e-07 AD=2.75125e-14 AS=2.6625e-14 PD=6.65e-07 PS=6.55e-07 $X=-13305 $Y=10720 $D=0
.ENDS
***************************************
.SUBCKT FA_2017 B A VDD GND Sum Cout Cin
** N=14 EP=7 IP=26 FDC=18
M0 6 B GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-11165 $Y=4275 $D=1
M1 5 A GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-11165 $Y=8455 $D=1
M2 10 8 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-3110 $Y=4275 $D=1
M3 11 9 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-3110 $Y=8455 $D=1
M4 Sum 10 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-2340 $Y=4275 $D=1
M5 Cout 11 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=-2340 $Y=8455 $D=1
M6 6 B VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-11165 $Y=5645 $D=0
M7 5 A VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-11165 $Y=9840 $D=0
M8 10 8 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-3110 $Y=5645 $D=0
M9 11 9 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-3110 $Y=9840 $D=0
M10 Sum 10 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-2340 $Y=5645 $D=0
M11 Cout 11 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=-2340 $Y=9840 $D=0
X20 GND VDD Cin 6 B 7 pass_mux $T=3830 -900 0 0 $X=-10350 $Y=8180
X21 GND VDD 7 A B 9 pass_mux $T=7750 -900 0 0 $X=-6430 $Y=8180
X22 GND VDD 7 5 A 8 pass_mux $T=7770 -5095 0 0 $X=-6410 $Y=3985
.ENDS
***************************************
