* SPICE NETLIST
***************************************

.SUBCKT PTAP_CDNS_593088949680
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NTAP_CDNS_593088949683
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TGFA_2010 B 2 A 4 Cout 6 Cin 8
** N=13 EP=8 IP=2 FDC=14
M0 13 A 9 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.655e-14 AS=1.62e-14 PD=7.7e-07 PS=5.4e-07 $X=-13995 $Y=4260 $D=1
M1 4 B 13 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.755e-14 AS=2.655e-14 PD=5.7e-07 PS=7.7e-07 $X=-13305 $Y=4260 $D=1
M2 Cout 10 A 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6875e-14 PD=5.45e-07 PS=5.55e-07 $X=-13270 $Y=3575 $D=1
M3 8 10 Cin 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6875e-14 PD=5.45e-07 PS=5.55e-07 $X=-12085 $Y=3570 $D=1
M4 10 9 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.125e-14 AS=1.1025e-14 PD=4.3e-07 PS=4.25e-07 $X=-11620 $Y=4290 $D=1
M5 Cout 9 Cin 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.665e-14 AS=1.665e-14 PD=5.5e-07 PS=5.5e-07 $X=-10755 $Y=3570 $D=1
M6 8 Cin 10 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.6425e-14 AS=1.6425e-14 PD=5.45e-07 PS=5.45e-07 $X=-10625 $Y=4280 $D=1
M7 9 A B 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.31e-14 AS=3.195e-14 PD=9.5e-07 PS=7.15e-07 $X=-13995 $Y=5790 $D=0
M8 A B 9 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.51e-14 AS=5.31e-14 PD=7.5e-07 PS=9.5e-07 $X=-13305 $Y=5790 $D=0
M9 Cout 9 A 2 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.375e-14 PD=7.05e-07 PS=7.35e-07 $X=-13260 $Y=1850 $D=0
M10 8 9 Cin 2 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.195e-14 AS=3.465e-14 PD=7.15e-07 PS=7.45e-07 $X=-12075 $Y=1850 $D=0
M11 10 9 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.205e-14 AS=2.16e-14 PD=6.05e-07 PS=6e-07 $X=-11620 $Y=5790 $D=0
M12 Cout 10 Cin 2 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.375e-14 PD=7.05e-07 PS=7.35e-07 $X=-10740 $Y=1850 $D=0
M13 8 Cin 9 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.465e-14 AS=3.06e-14 PD=7.45e-07 PS=7e-07 $X=-10625 $Y=5790 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=13 EP=13 IP=16 FDC=28
X0 3 13 4 11 5 12 6 1 TGFA_2010 $T=0 0 0 0 $X=-15460 $Y=1610
X1 7 13 8 11 9 12 10 2 TGFA_2010 $T=6000 0 0 0 $X=-9460 $Y=1610
.ENDS
***************************************
.SUBCKT and2 B GND VDD Y
** N=7 EP=4 IP=0 FDC=6
M0 7 A GND GND NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.88e-14 PD=6.4e-07 PS=6.8e-07 $X=3340 $Y=6545 $D=1
M1 6 B 7 GND NMOS_VTL L=5e-08 W=1.8e-07 AD=3.06e-14 AS=2.52e-14 PD=7e-07 PS=6.4e-07 $X=3720 $Y=6545 $D=1
M2 Y 6 GND GND NMOS_VTL L=5.25e-08 W=9e-08 AD=1.1475e-14 AS=1.2375e-14 PD=4.35e-07 PS=4.55e-07 $X=5155 $Y=6635 $D=1
M3 6 A VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=4.41e-14 AS=2.88e-14 PD=8.5e-07 PS=6.8e-07 $X=3340 $Y=7995 $D=0
M4 VDD B 6 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=3.555e-14 AS=4.41e-14 PD=7.55e-07 PS=8.5e-07 $X=3930 $Y=7995 $D=0
M5 Y 6 VDD VDD PMOS_VTL L=5.25e-08 W=1.8e-07 AD=2.295e-14 AS=2.025e-14 PD=6.15e-07 PS=5.85e-07 $X=5155 $Y=8005 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=8 FDC=12
X0 1 2 3 4 and2 $T=0 12280 1 0 $X=2840 $Y=3650
X1 5 6 7 8 and2 $T=0 0 0 0 $X=2840 $Y=6250
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=8 FDC=12
X0 1 2 3 4 and2 $T=0 0 0 0 $X=2840 $Y=6250
X1 5 6 7 8 and2 $T=3000 0 0 0 $X=5840 $Y=6250
.ENDS
***************************************
.SUBCKT W_Mul GND X1 Y0 Y3 Y2 Y1 P7 P0 P1 P2 P4 P5 P6 P3 VDD
** N=57 EP=15 IP=152 FDC=264
X4 9 VDD 11 GND 24 VDD 9 16 TGFA_2010 $T=37790 21405 1 0 $X=22330 $Y=15015
X5 7 47 10 GND 18 VDD 8 17 TGFA_2010 $T=37790 26185 1 0 $X=22330 $Y=19795
X6 30 VDD 32 GND 53 VDD GND P3 TGFA_2010 $T=52790 11845 1 0 $X=37330 $Y=5455
X7 28 VDD 26 GND 54 VDD 53 P4 TGFA_2010 $T=52790 16625 1 0 $X=37330 $Y=10235
X8 P1 P2 12 15 23 GND 23 25 30 GND GND VDD VDD ICV_1 $T=40790 11845 1 0 $X=25330 $Y=5455
X9 25 32 13 GND 52 14 16 19 28 52 GND VDD VDD ICV_1 $T=40790 16625 1 0 $X=25330 $Y=10235
X10 26 P5 24 17 29 GND 29 27 55 54 GND VDD VDD ICV_1 $T=46790 21405 1 0 $X=31330 $Y=15015
X11 27 P6 21 22 31 18 31 20 P7 55 GND VDD 57 ICV_1 $T=46790 26185 1 0 $X=31330 $Y=19795
X12 Y3 X1 43 10 Y0 GND 44 9 ICV_2 $T=16420 23545 1 0 $X=19260 $Y=14915
X13 Y1 GND 45 8 Y2 GND 43 7 ICV_2 $T=16420 28325 1 0 $X=19260 $Y=19695
X14 Y3 GND VDD 20 Y3 GND VDD 19 ICV_2 $T=25420 23545 1 0 $X=28260 $Y=14915
X15 Y2 GND 47 21 Y3 GND VDD 22 ICV_2 $T=25420 28325 1 0 $X=28260 $Y=19695
X16 Y0 GND P0 P0 Y1 GND 48 15 ICV_3 $T=16420 13985 1 0 $X=19260 $Y=5355
X17 Y2 GND 49 GND Y0 X1 50 12 ICV_3 $T=16420 1705 0 0 $X=19260 $Y=7955
X18 Y2 X1 49 11 Y1 X1 50 13 ICV_3 $T=16420 18765 1 0 $X=19260 $Y=10135
X19 Y1 GND 44 9 Y0 GND 51 14 ICV_3 $T=16420 6485 0 0 $X=19260 $Y=12735
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
